library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity IM is
    port(
        CLK : in std_logic;
        IMA : in std_logic_vector(31 downto 0);
        IMOut : out std_logic_vector(31 downto 0)
    );
end IM;

architecture RTL of IM is

begin
                  -- R Type : < op ><rs ><rt ><rd ><sha><func>
                  -- I Type : < op ><rs ><rt ><   imm/addr   >
                  -- J Type : < op ><          addr          >
    IMo : process(IMA(7 downto 2))
    begin
        case (IMA(7 downto 2)) is
            when "000000" => 
                IMOut <= "00000111101111011111111111111100";
            when "000001" => 
                IMOut <= "00001111101111110000000000000000";
            when "000010" => 
                IMOut <= "00000100000111100000000000001000";
            when "000011" => 
                IMOut <= "00011000000000000000000000001000";
            when "000100" => 
                IMOut <= "00000100010111100000000000000000";
            when "000101" => 
                IMOut <= "00001011101111110000000000000000";
            when "000110" => 
                IMOut <= "00000111101111010000000000000100";
            when "000111" => 
                IMOut <= "00011111111000000000000000000000";
            when "001000" => 
                IMOut <= "00010011110000000000000000001111";
            when "001001" => 
                IMOut <= "00000111101111011111111111111000";
            when "001010" => 
                IMOut <= "00001111101111110000000000000100";
            when "001011" => 
                IMOut <= "00001111101111100000000000000000";
            when "001100" => 
                IMOut <= "00000111110111101111111111111111";
            when "001101" => 
                IMOut <= "00011000000000000000000000001000";
            when "001110" => 
                IMOut <= "00001011101111110000000000000100";
            when "001111" => 
                IMOut <= "00001011101111100000000000000000";
            when "010000" => 
                IMOut <= "00000111101111010000000000001000";
            when "010001" => 
                IMOut <= "00000100000000110000000000000000";
            when "010010" => 
                IMOut <= "00000000011000100001100000000000";
            when "010011" => 
                IMOut <= "00000111110111101111111111111111";
            when "010100" => 
                IMOut <= "00010011110000000000000000000001";
            when "010101" => 
                IMOut <= "00010100000000000000000000010010";
            when "010110" => 
                IMOut <= "00000100011000100000000000000000";
            when "010111" => 
                IMOut <= "00011111111000000000000000000000";
            when "011000" => 
                IMOut <= "00000100000000100000000000000001";
            when "011001" => 
                IMOut <= "00011111111000000000000000000000";

            when others =>  -- nop : add $0,$0,$0
                    IMOut <= "00000000000000000000000000000000";
        end case;
    end process;

end RTL;
